`define NRSPACES 14
`define PER_RSP [`NRSPACES-1:0]
`define BITNESS 64
`define WORD [`BITNESS-1:0]
